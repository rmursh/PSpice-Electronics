Inverting Amplifier
**CIRCUIT DESCRIPTION**
*POWER SUPPLY*
Vin 5 0 SIN(0 100m 1k 0 0)

*ELEMENTS*
R1 0 2 5K
R2 5 1 5K
R3 2 6 100K
RL 6 0 1K
X1 1 2 3 OPAMP
D1 3 6 dmodel

.model dmodel d(Is=1e-9 n=1.8)


**ANALYSIS REQUUEST**
.TRAN 1u 5m 0 1u

**OUTPUT REQUEST**
.PLOT TRAN V(1,0), V(6,0)
.PROBE


*             non-inverting input
*             | inverting input
*             | | output
*             | | |
.SUBCKT OPAMP 1 2 3


*CIRCUIT DESCRIPTION

*SOURCE
EV3 4 0 1 2 10K
Rin 1 2 1MEG
Rout 4 3 50


.ENDS OPAMP




.END