*CASCODE AMPLIFIER*
Vdd 5 0 DC 15
*Vtst 1 0 ac 1m 0
Vsig 1 0 sin 0 0.00 50K 0 0

*RESISTOR ELEMENTS*
Rsig 1 2 1K 
R1 3 0 180K
R2 4 3 56K 
R3 5 4 270K 
RC 5 6 3.9K 
RE 8 0 3.3K 
RL 9 0 1K 

*CAPACITOR ELEMENTS*
C1 3 2 3.3u 
CB 4 0 4.7u  
C2 9 6 3.3u 
CE 8 0 100u 

*BJT*
Q1 7 3 8 QMPS2222A
Q2 6 4 7 QMPS2222A


*MODEL SPECIFICATION*
*MPS2222A MCE 1/26/96
*Si 625mW 40V 600mA 300MHz pkg:TO-92 1,2,3
.MODEL QMPS2222A NPN (IS=.504F NF=1 BF=339 VAF=113 IKF=.36 ISE=1.63P NE=2
+ BR=4 NR=1 VAR=24 IKR=.54 RE=.173 RB=.692 RC=69.2M XTB=1.5
+ CJE=23.5P VJE=1.1 MJE=.5 CJC=10.6P VJC=.3 MJC=.3 TF=521P TR=272N)

*ANALYSIS REQUEST*

.op
*.ac dec 10 1  10G	
.tran 1n 0.1m

*OUTPUT REQUEST*
.probe  

.end