Question 1 part a
*Plot Vsig, Vi, Vo, Io

*Source
VSigV 1 0 SIN(0 1 10)

*circuit description
RSigR 2 1 50
CCap1 3 2 1uF
RRes1 3 0 100k
RRes2 3 0 100k


GmVi 4 0 3 0 50m
RResD 4 0 10k
CCap2 5 4 1uF
RResL 5 0 10k


*analysis request
.TRAN 1m 1 0 1m

.PLOT TRAN V(1,0) V(5,0)
.PROBE

.END