Operational Amplifier Model
**	CIRCUIT DESCRIPTION**
*POWER SUPPLY*
Vin-diff 6 0 SIN(0 5m 1k 0 0)
Vcm 5 0 1
EV1 1 5 6 0 0.5
EV2 5 2 6 0 0.5



*ELEMENTS*
X1 1 2 3 OPAMP
RL 3 0 1K
R1 6 0 1K


**ANALYSIS REQUESTS**
.TRAN 1u 1m 0 1u

**OUTPUT REQUEST**
.PLOT TRAN V(1,0) V(6,0)
.PROBE



*             non-inverting input
*             | inverting input
*             | | output
*             | | |
.SUBCKT OPAMP 1 2 3


*CIRCUIT DESCRIPTION

*SOURCE
EV3 4 0 1 2 10K
Rin 1 2 1MEG
Rout 4 3 50


.ENDS OPAMP

.END