Biasing MOSFET Amplifier
**CIRCUIT DESCRIPTION**
*VOLTAGE SUPPLY*
VDD 2 0 DC 20
Vsig 8 0 AC 5m 0

*RESISTOR ELEMENTS*
Rsig 8 7 50
R1 1 0 10MEG
R2 2 1 10MEG 
RD1 4 0 2.5K
RS1 2 3 1K
RS2 6 0 500
RD2 2 5 1K
RL 9 0 1K

*CAPACITORS*

C1 7 1 100u
C2 9 5 100u
CS1 2 3 100u
CS2 6 0 100u 



*MOS*
M1 4 1 3 3 PFET L=20u W=350u

M2 5 4 6 6 NFET L=20u W=100u

.MODEL nfet NMOS LEVEL=3 PHI=0.600000 TOX=2.1200E-08
+ XJ=0.200000U TPG=1 VTO=0.7860 DELTA=6.9670E-01
+ LD=1.6470E-07 KP=9.6379E-05 UO=591.7 THETA=8.1220E-02
+ RSH=8.5450E+01 GAMMA=0.5863 NSUB=1.6160E+16
+ NFS=5.0000E+12 VMAX=2.0820E+05 ETA=7.0660E-02
+ KAPPA=1.3960E-01 CGDO=4.0241E-10 CGSO=4.0241E-10
+ CGBO=3.6144E-10 CJ=3.8541E-04 MJ=1.1854
+ CJSW=1.3940E-10 MJSW=0.125195 PB=0.800000

.MODEL pfet PMOS LEVEL=3 PHI=0.600000 TOX=2.1200E-08
+ XJ=0.200000U TPG=-1 VTO=-0.9056 DELTA=1.5200E+00
+ LD=2.2000E-08 KP=2.9352E-05 UO=180.2 THETA=1.2480E-01
+ RSH=1.0470E+02 GAMMA=0.4863 NSUB=1.8900E+16
+ NFS=3.46E+12 VMAX=3.7320E+05 ETA=1.6410E-01
+ KAPPA=9.6940E+00 CGDO=5.3752E-11 CGSO=5.3752E-11
+ CGBO=3.3650E-10 CJ=4.8447E-04 MJ=0.5027
+ CJSW=1.6457E-10 MJSW=0.217168 PB=0.850000


*ANALYSIS REQUEST*
.AC DEC 10 1m 1G

*OUTPUT REQUEST*

.PROBE

.END